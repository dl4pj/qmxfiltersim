.title QMX FILTER SIMULATION
* .include "qmxfilters.lib"

* SWEEP:


.control
set hcopydevtype=svg

set start = 1Meg
set stop = 150Meg
set points = 10000

foreach dut bpf6m bpf10m bpf15m bpf20m lpf6m lpf10m lpf15m lpf20m lpfbpf6m lpfbpf10m lpfbpf15m lpfbpf20m

circbyline QMX Filters
circbyline .include "qmxfilters.lib"
circbyline V1  p1 0 DC 0 AC 1 portnum 1
circbyline V2  p2 0 DC 0      portnum 2
circbyline X1 p1 p2 $dut

circbyline .end
sp lin $points $start $stop
set filename={$dut}.svg
let vswr = ( 1+ abs(s_1_1) ) / (1.000000001 - abs(s_1_1)) 
hardcopy ./out/$filename vdb(s_1_1) vdb(s_2_1) vswr ylimit -120 20 xlabel 'Frequency' ylabel 'Magnitude in dB / VSWR' title $dut
remcirc
reset

end ; foreach


.endc
.end